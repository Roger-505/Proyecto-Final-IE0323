/* Red iterativa 
   -------------
    Conductual */

module redIterativa 
#( parameter N = 3 ) 
(
    input [N-1:0]A, [N-1:0]B 
);
    
endmodule