/* Definición de módulo para la celda típica de la 
   red iterativa analizando las palabras de derecha 
   a izquierda*/

module celdaTipica (
    input p, Ai, Bi,
    output P
); 
always @(p or Ai or Bi)
begin
    

end 
endendmodule